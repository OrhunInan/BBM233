`timescale 1ns/10ps

module multiplier_tb;

reg [2:0] A, B;
wire [5:0] Out;

multiplier UUT(.A(A), .B(B), .P(Out));

initial begin
    
    $dumpfile("multiplier.vcd");
	$dumpvars;

    A = 000; B = 000;
    #10; A = 000; B = 001;
    #10; A = 000; B = 010;
    #10; A = 000; B = 011;
    #10; A = 000; B = 100;
    #10; A = 000; B = 101;
    #10; A = 000; B = 110;
    #10; A = 000; B = 111;
	#10; A = 001; B = 000;
	#10; A = 001; B = 001;
    #10; A = 001; B = 010;
    #10; A = 001; B = 011;
    #10; A = 001; B = 100;
    #10; A = 001; B = 101;
    #10; A = 001; B = 110;
    #10; A = 001; B = 111;
	#10; A = 010; B = 000;
	#10; A = 010; B = 001;
    #10; A = 010; B = 010;
    #10; A = 010; B = 011;
    #10; A = 010; B = 100;
    #10; A = 010; B = 101;
    #10; A = 010; B = 110;
    #10; A = 010; B = 111;
	#10; A = 011; B = 000;
	#10; A = 011; B = 001;
    #10; A = 011; B = 010;
    #10; A = 011; B = 011;
    #10; A = 011; B = 100;
    #10; A = 011; B = 101;
    #10; A = 011; B = 110;
    #10; A = 011; B = 111;
	#10; A = 100; B = 000;
	#10; A = 100; B = 001;
    #10; A = 100; B = 010;
    #10; A = 100; B = 011;
    #10; A = 100; B = 100;
    #10; A = 100; B = 101;
    #10; A = 100; B = 110;
    #10; A = 100; B = 111;
	#10; A = 101; B = 000;
	#10; A = 101; B = 001;
    #10; A = 101; B = 010;
    #10; A = 101; B = 011;
    #10; A = 101; B = 100;
    #10; A = 101; B = 101;
    #10; A = 101; B = 110;
    #10; A = 101; B = 111;
	#10; A = 110; B = 000;
	#10; A = 110; B = 001;
    #10; A = 110; B = 010;
    #10; A = 110; B = 011;
    #10; A = 110; B = 100;
    #10; A = 110; B = 101;
    #10; A = 110; B = 110;
    #10; A = 110; B = 111;
	#10; A = 111; B = 000;
	#10; A = 111; B = 001;
    #10; A = 111; B = 010;
    #10; A = 111; B = 011;
    #10; A = 111; B = 100;
    #10; A = 111; B = 101;
    #10; A = 111; B = 110;
    #10; A = 111; B = 111;
    #10; $finish;
end

endmodule
